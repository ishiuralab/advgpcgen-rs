module testbench();
    reg [6:0] src0;
    reg [3:0] src2;
    reg [0:0] src3;
    wire [4:0] dst;
    wire [4:0] exp;
    wire test;
    gpc1407_5 gpc1407_5(
        .src0(src0),
        .src2(src2),
        .src3(src3),
        .dst(dst)
    );
    assign exp = src0[0] * 1 + src0[1] * 1 + src0[2] * 1 + src0[3] * 1 + src0[4] * 1 + src0[5] * 1 + src0[6] * 1 + src2[0] * 4 + src2[1] * 4 + src2[2] * 4 + src2[3] * 4 + src3[0] * 8;
    assign test = dst == exp;
    initial begin
        $monitor("src0:0x%x, src2:0x%x, src3:0x%x, dst:0x%x, exp:0x%x, test:%x", src0, src2, src3, dst, exp, test);
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h100;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h101;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h102;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h103;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h104;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h105;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h106;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h107;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h108;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h109;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h10f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h110;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h111;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h112;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h113;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h114;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h115;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h116;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h117;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h118;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h119;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h11f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h120;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h121;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h122;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h123;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h124;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h125;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h126;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h127;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h128;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h129;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h12f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h130;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h131;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h132;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h133;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h134;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h135;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h136;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h137;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h138;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h139;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h13f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h140;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h141;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h142;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h143;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h144;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h145;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h146;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h147;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h148;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h149;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h14f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h150;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h151;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h152;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h153;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h154;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h155;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h156;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h157;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h158;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h159;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h15f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h160;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h161;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h162;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h163;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h164;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h165;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h166;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h167;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h168;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h169;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h16f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h170;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h171;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h172;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h173;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h174;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h175;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h176;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h177;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h178;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h179;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h17f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h180;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h181;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h182;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h183;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h184;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h185;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h186;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h187;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h188;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h189;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h18f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h190;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h191;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h192;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h193;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h194;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h195;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h196;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h197;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h198;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h199;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h19f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h1ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h200;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h201;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h202;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h203;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h204;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h205;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h206;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h207;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h208;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h209;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h20f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h210;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h211;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h212;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h213;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h214;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h215;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h216;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h217;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h218;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h219;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h21f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h220;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h221;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h222;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h223;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h224;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h225;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h226;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h227;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h228;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h229;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h22f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h230;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h231;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h232;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h233;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h234;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h235;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h236;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h237;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h238;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h239;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h23f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h240;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h241;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h242;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h243;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h244;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h245;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h246;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h247;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h248;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h249;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h24f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h250;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h251;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h252;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h253;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h254;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h255;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h256;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h257;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h258;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h259;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h25f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h260;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h261;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h262;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h263;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h264;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h265;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h266;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h267;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h268;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h269;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h26f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h270;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h271;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h272;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h273;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h274;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h275;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h276;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h277;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h278;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h279;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h27f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h280;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h281;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h282;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h283;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h284;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h285;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h286;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h287;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h288;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h289;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h28f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h290;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h291;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h292;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h293;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h294;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h295;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h296;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h297;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h298;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h299;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h29f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h2ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h300;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h301;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h302;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h303;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h304;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h305;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h306;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h307;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h308;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h309;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h30f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h310;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h311;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h312;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h313;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h314;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h315;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h316;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h317;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h318;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h319;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h31f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h320;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h321;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h322;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h323;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h324;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h325;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h326;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h327;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h328;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h329;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h32f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h330;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h331;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h332;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h333;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h334;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h335;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h336;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h337;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h338;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h339;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h33f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h340;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h341;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h342;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h343;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h344;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h345;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h346;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h347;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h348;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h349;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h34f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h350;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h351;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h352;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h353;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h354;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h355;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h356;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h357;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h358;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h359;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h35f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h360;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h361;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h362;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h363;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h364;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h365;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h366;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h367;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h368;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h369;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h36f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h370;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h371;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h372;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h373;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h374;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h375;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h376;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h377;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h378;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h379;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h37f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h380;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h381;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h382;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h383;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h384;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h385;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h386;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h387;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h388;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h389;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h38f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h390;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h391;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h392;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h393;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h394;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h395;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h396;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h397;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h398;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h399;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h39f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h3ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h400;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h401;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h402;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h403;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h404;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h405;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h406;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h407;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h408;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h409;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h40f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h410;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h411;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h412;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h413;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h414;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h415;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h416;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h417;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h418;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h419;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h41f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h420;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h421;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h422;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h423;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h424;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h425;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h426;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h427;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h428;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h429;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h42f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h430;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h431;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h432;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h433;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h434;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h435;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h436;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h437;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h438;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h439;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h43f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h440;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h441;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h442;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h443;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h444;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h445;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h446;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h447;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h448;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h449;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h44f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h450;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h451;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h452;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h453;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h454;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h455;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h456;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h457;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h458;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h459;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h45f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h460;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h461;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h462;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h463;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h464;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h465;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h466;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h467;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h468;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h469;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h46f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h470;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h471;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h472;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h473;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h474;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h475;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h476;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h477;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h478;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h479;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h47f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h480;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h481;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h482;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h483;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h484;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h485;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h486;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h487;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h488;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h489;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h48f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h490;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h491;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h492;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h493;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h494;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h495;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h496;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h497;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h498;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h499;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h49f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h4ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h500;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h501;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h502;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h503;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h504;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h505;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h506;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h507;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h508;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h509;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h50f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h510;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h511;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h512;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h513;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h514;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h515;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h516;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h517;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h518;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h519;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h51f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h520;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h521;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h522;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h523;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h524;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h525;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h526;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h527;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h528;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h529;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h52f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h530;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h531;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h532;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h533;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h534;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h535;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h536;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h537;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h538;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h539;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h53f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h540;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h541;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h542;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h543;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h544;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h545;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h546;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h547;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h548;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h549;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h54f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h550;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h551;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h552;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h553;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h554;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h555;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h556;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h557;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h558;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h559;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h55f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h560;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h561;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h562;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h563;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h564;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h565;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h566;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h567;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h568;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h569;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h56f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h570;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h571;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h572;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h573;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h574;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h575;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h576;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h577;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h578;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h579;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h57f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h580;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h581;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h582;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h583;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h584;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h585;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h586;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h587;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h588;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h589;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h58f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h590;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h591;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h592;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h593;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h594;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h595;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h596;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h597;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h598;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h599;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h59f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h5ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h600;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h601;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h602;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h603;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h604;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h605;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h606;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h607;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h608;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h609;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h60f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h610;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h611;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h612;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h613;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h614;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h615;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h616;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h617;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h618;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h619;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h61f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h620;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h621;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h622;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h623;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h624;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h625;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h626;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h627;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h628;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h629;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h62f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h630;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h631;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h632;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h633;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h634;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h635;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h636;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h637;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h638;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h639;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h63f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h640;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h641;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h642;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h643;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h644;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h645;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h646;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h647;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h648;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h649;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h64f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h650;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h651;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h652;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h653;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h654;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h655;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h656;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h657;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h658;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h659;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h65f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h660;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h661;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h662;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h663;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h664;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h665;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h666;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h667;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h668;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h669;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h66f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h670;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h671;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h672;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h673;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h674;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h675;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h676;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h677;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h678;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h679;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h67f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h680;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h681;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h682;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h683;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h684;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h685;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h686;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h687;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h688;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h689;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h68f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h690;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h691;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h692;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h693;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h694;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h695;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h696;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h697;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h698;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h699;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h69f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h6ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h700;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h701;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h702;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h703;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h704;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h705;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h706;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h707;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h708;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h709;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h70f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h710;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h711;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h712;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h713;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h714;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h715;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h716;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h717;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h718;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h719;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h71f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h720;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h721;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h722;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h723;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h724;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h725;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h726;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h727;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h728;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h729;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h72f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h730;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h731;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h732;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h733;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h734;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h735;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h736;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h737;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h738;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h739;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h73f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h740;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h741;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h742;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h743;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h744;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h745;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h746;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h747;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h748;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h749;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h74f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h750;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h751;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h752;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h753;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h754;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h755;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h756;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h757;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h758;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h759;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h75f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h760;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h761;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h762;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h763;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h764;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h765;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h766;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h767;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h768;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h769;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h76f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h770;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h771;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h772;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h773;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h774;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h775;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h776;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h777;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h778;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h779;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h77f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h780;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h781;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h782;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h783;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h784;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h785;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h786;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h787;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h788;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h789;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h78f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h790;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h791;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h792;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h793;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h794;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h795;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h796;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h797;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h798;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h799;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h79f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h7ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h800;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h801;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h802;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h803;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h804;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h805;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h806;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h807;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h808;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h809;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h80f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h810;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h811;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h812;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h813;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h814;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h815;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h816;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h817;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h818;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h819;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h81f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h820;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h821;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h822;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h823;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h824;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h825;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h826;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h827;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h828;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h829;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h82f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h830;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h831;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h832;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h833;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h834;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h835;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h836;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h837;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h838;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h839;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h83f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h840;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h841;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h842;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h843;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h844;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h845;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h846;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h847;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h848;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h849;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h84f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h850;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h851;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h852;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h853;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h854;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h855;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h856;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h857;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h858;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h859;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h85f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h860;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h861;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h862;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h863;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h864;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h865;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h866;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h867;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h868;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h869;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h86f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h870;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h871;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h872;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h873;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h874;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h875;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h876;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h877;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h878;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h879;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h87f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h880;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h881;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h882;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h883;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h884;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h885;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h886;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h887;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h888;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h889;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h88f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h890;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h891;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h892;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h893;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h894;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h895;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h896;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h897;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h898;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h899;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h89f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h8ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h900;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h901;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h902;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h903;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h904;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h905;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h906;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h907;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h908;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h909;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h90f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h910;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h911;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h912;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h913;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h914;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h915;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h916;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h917;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h918;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h919;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h91f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h920;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h921;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h922;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h923;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h924;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h925;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h926;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h927;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h928;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h929;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h92f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h930;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h931;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h932;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h933;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h934;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h935;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h936;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h937;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h938;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h939;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h93f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h940;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h941;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h942;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h943;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h944;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h945;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h946;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h947;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h948;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h949;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h94f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h950;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h951;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h952;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h953;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h954;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h955;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h956;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h957;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h958;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h959;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h95f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h960;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h961;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h962;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h963;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h964;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h965;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h966;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h967;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h968;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h969;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h96f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h970;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h971;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h972;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h973;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h974;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h975;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h976;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h977;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h978;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h979;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h97f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h980;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h981;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h982;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h983;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h984;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h985;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h986;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h987;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h988;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h989;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h98f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h990;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h991;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h992;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h993;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h994;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h995;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h996;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h997;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h998;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h999;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h99f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'h9ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha00;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha01;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha02;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha03;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha04;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha05;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha06;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha07;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha08;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha09;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha0f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'ha9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haa9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haaa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haaf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hab9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'habb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'habc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'habd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'habe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'habf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hac9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hacb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hacc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hacd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hace;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hacf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'had9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hada;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hadb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hadc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hadd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hade;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hadf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hae9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haeb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haf9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hafa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hafb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hafc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hafd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hafe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'haff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb00;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb01;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb02;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb03;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb04;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb05;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb06;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb07;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb08;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb09;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb0f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hb9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hba9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbaa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbaf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbbb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbbc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbbd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbbe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbbf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbc9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbcb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbcc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbcd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbcf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbd9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbdb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbdc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbdd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbde;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbdf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbe9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbeb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbf9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbfa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbfb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbfc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbfd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbfe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hbff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc00;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc01;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc02;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc03;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc04;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc05;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc06;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc07;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc08;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc09;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc0f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hc9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hca9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcaa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcaf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcbb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcbc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcbd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcbe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcbf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcc9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hccb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hccc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hccd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hccf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcd9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcdb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcdc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcdd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcde;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcdf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hce9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hceb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hced;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcf9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcfa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcfb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcfc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcfd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcfe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hcff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd00;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd01;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd02;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd03;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd04;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd05;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd06;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd07;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd08;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd09;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd0f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hd9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hda9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdaa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdaf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdbb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdbc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdbd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdbe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdbf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdc9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdcb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdcc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdcd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdcf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdd9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hddb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hddc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hddd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdde;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hddf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hde9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdeb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hded;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdf9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdfa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdfb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdfc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdfd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdfe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hdff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he00;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he01;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he02;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he03;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he04;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he05;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he06;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he07;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he08;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he09;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he0f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'he9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hea9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heaa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'head;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heaf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hebb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hebc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hebd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hebe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hebf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hec9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hecb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hecc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hecd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hece;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hecf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hed9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hedb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hedc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hedd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hede;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hedf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hee9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heeb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hef9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hefa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hefb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hefc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hefd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hefe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'heff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf00;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf01;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf02;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf03;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf04;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf05;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf06;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf07;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf08;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf09;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf0f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hf9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfa9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfaa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfaf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfbb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfbc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfbd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfbe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfbf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfc9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfcb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfcc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfcd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfcf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfd9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfdb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfdc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfdd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfde;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfdf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfe9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfeb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hff9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hffa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hffb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hffc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hffd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hffe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 12'hfff;
        #1
        $finish();
    end
endmodule
