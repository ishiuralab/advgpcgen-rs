module testbench();
    reg [0:0] src0;
    reg [6:0] src1;
    reg [1:0] src3;
    wire [4:0] dst;
    wire [4:0] exp;
    wire test;
    gpc2071_5 gpc2071_5(
        .src0(src0),
        .src1(src1),
        .src3(src3),
        .dst(dst)
    );
    assign exp = src0[0] * 1 + src1[0] * 2 + src1[1] * 2 + src1[2] * 2 + src1[3] * 2 + src1[4] * 2 + src1[5] * 2 + src1[6] * 2 + src3[0] * 8 + src3[1] * 8;
    assign test = dst == exp;
    initial begin
        $monitor("src0:0x%x, src1:0x%x, src3:0x%x, dst:0x%x, exp:0x%x, test:%x", src0, src1, src3, dst, exp, test);
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h40;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h41;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h42;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h43;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h44;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h45;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h46;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h47;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h48;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h49;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h4f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h50;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h51;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h52;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h53;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h54;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h55;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h56;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h57;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h58;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h59;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h5f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h60;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h61;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h62;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h63;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h64;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h65;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h66;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h67;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h68;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h69;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h6f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h70;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h71;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h72;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h73;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h74;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h75;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h76;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h77;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h78;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h79;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h7f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h80;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h81;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h82;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h83;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h84;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h85;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h86;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h87;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h88;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h89;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h8f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h90;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h91;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h92;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h93;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h94;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h95;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h96;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h97;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h98;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h99;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h9f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'ha9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'haa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hab;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hac;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'had;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hae;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'haf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hb9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hba;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hbb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hbc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hbd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hbe;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hbf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hc9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hca;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hcb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hcc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hcd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hce;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hcf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hd9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hda;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hdb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hdc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hdd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hde;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hdf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'he9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hea;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'heb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hec;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hed;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hee;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hef;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hf9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hfa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hfb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hfc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hfd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hfe;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'hff;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h100;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h101;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h102;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h103;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h104;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h105;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h106;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h107;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h108;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h109;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h10f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h110;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h111;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h112;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h113;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h114;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h115;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h116;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h117;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h118;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h119;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h11f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h120;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h121;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h122;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h123;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h124;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h125;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h126;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h127;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h128;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h129;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h12f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h130;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h131;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h132;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h133;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h134;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h135;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h136;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h137;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h138;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h139;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h13f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h140;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h141;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h142;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h143;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h144;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h145;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h146;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h147;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h148;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h149;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h14f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h150;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h151;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h152;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h153;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h154;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h155;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h156;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h157;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h158;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h159;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h15f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h160;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h161;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h162;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h163;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h164;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h165;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h166;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h167;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h168;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h169;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h16f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h170;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h171;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h172;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h173;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h174;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h175;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h176;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h177;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h178;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h179;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h17f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h180;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h181;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h182;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h183;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h184;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h185;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h186;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h187;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h188;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h189;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h18f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h190;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h191;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h192;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h193;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h194;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h195;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h196;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h197;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h198;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h199;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h19f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1a9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1aa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ab;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ac;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ad;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ae;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1af;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1b9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ba;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1bb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1bc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1bd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1be;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1bf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1c9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ca;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1cb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1cc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1cd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ce;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1cf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1d9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1da;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1db;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1dc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1dd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1de;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1df;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1e9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ea;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1eb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ec;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ed;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ee;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ef;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1f9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1fa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1fb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1fc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1fd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1fe;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h1ff;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h200;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h201;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h202;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h203;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h204;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h205;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h206;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h207;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h208;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h209;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h20f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h210;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h211;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h212;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h213;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h214;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h215;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h216;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h217;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h218;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h219;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h21f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h220;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h221;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h222;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h223;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h224;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h225;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h226;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h227;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h228;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h229;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h22f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h230;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h231;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h232;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h233;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h234;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h235;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h236;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h237;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h238;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h239;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h23f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h240;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h241;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h242;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h243;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h244;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h245;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h246;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h247;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h248;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h249;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h24f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h250;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h251;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h252;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h253;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h254;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h255;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h256;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h257;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h258;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h259;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h25f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h260;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h261;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h262;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h263;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h264;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h265;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h266;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h267;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h268;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h269;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h26f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h270;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h271;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h272;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h273;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h274;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h275;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h276;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h277;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h278;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h279;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h27f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h280;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h281;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h282;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h283;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h284;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h285;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h286;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h287;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h288;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h289;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h28f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h290;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h291;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h292;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h293;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h294;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h295;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h296;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h297;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h298;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h299;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h29f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2a9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2aa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ab;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ac;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ad;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ae;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2af;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2b9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ba;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2bb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2bc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2bd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2be;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2bf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2c9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ca;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2cb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2cc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2cd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ce;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2cf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2d9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2da;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2db;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2dc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2dd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2de;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2df;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2e9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ea;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2eb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ec;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ed;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ee;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ef;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2f9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2fa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2fb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2fc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2fd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2fe;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h2ff;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h300;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h301;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h302;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h303;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h304;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h305;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h306;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h307;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h308;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h309;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h30f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h310;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h311;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h312;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h313;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h314;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h315;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h316;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h317;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h318;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h319;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h31f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h320;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h321;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h322;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h323;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h324;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h325;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h326;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h327;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h328;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h329;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h32f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h330;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h331;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h332;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h333;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h334;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h335;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h336;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h337;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h338;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h339;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h33f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h340;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h341;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h342;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h343;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h344;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h345;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h346;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h347;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h348;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h349;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h34f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h350;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h351;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h352;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h353;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h354;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h355;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h356;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h357;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h358;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h359;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h35f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h360;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h361;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h362;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h363;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h364;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h365;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h366;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h367;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h368;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h369;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h36f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h370;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h371;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h372;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h373;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h374;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h375;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h376;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h377;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h378;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h379;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h37f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h380;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h381;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h382;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h383;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h384;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h385;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h386;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h387;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h388;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h389;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h38f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h390;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h391;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h392;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h393;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h394;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h395;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h396;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h397;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h398;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h399;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39a;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39b;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39c;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39d;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39e;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h39f;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3a9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3aa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ab;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ac;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ad;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ae;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3af;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3b9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ba;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3bb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3bc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3bd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3be;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3bf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3c9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ca;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3cb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3cc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3cd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ce;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3cf;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3d9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3da;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3db;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3dc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3dd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3de;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3df;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3e9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ea;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3eb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ec;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ed;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ee;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ef;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f0;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f1;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f2;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f3;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f4;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f5;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f6;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f7;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f8;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3f9;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3fa;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3fb;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3fc;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3fd;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3fe;
        #1
        {src3[1], src3[0], src1[6], src1[5], src1[4], src1[3], src1[2], src1[1], src1[0], src0[0]} <= 10'h3ff;
        #1
        $finish();
    end
endmodule
