module testbench();
    reg [5:0] src0;
    reg [3:0] src2;
    reg [0:0] src3;
    wire [4:0] dst;
    wire [4:0] exp;
    wire test;
    gpc1406_5 gpc1406_5(
        .src0(src0),
        .src2(src2),
        .src3(src3),
        .dst(dst)
    );
    assign exp = src0[0] * 1 + src0[1] * 1 + src0[2] * 1 + src0[3] * 1 + src0[4] * 1 + src0[5] * 1 + src2[0] * 4 + src2[1] * 4 + src2[2] * 4 + src2[3] * 4 + src3[0] * 8;
    assign test = dst == exp;
    initial begin
        $monitor("src0:0x%x, src2:0x%x, src3:0x%x, dst:0x%x, exp:0x%x, test:%x", src0, src2, src3, dst, exp, test);
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h80;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h81;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h82;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h83;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h84;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h85;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h86;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h87;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h88;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h89;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h8f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h90;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h91;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h92;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h93;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h94;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h95;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h96;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h97;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h98;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h99;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h9f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'ha9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'haa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'had;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'haf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hb9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hbb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hbc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hbd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hbe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hbf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hc9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hcb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hcc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hcd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hcf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hd9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hda;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hdb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hdc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hdd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hde;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hdf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'he9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'heb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hf9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hfa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hfb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hfc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hfd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hfe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'hff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h100;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h101;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h102;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h103;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h104;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h105;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h106;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h107;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h108;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h109;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h10f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h110;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h111;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h112;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h113;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h114;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h115;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h116;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h117;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h118;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h119;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h11f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h120;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h121;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h122;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h123;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h124;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h125;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h126;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h127;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h128;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h129;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h12f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h130;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h131;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h132;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h133;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h134;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h135;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h136;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h137;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h138;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h139;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h13f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h140;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h141;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h142;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h143;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h144;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h145;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h146;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h147;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h148;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h149;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h14f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h150;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h151;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h152;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h153;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h154;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h155;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h156;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h157;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h158;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h159;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h15f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h160;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h161;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h162;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h163;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h164;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h165;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h166;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h167;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h168;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h169;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h16f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h170;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h171;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h172;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h173;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h174;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h175;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h176;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h177;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h178;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h179;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h17f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h180;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h181;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h182;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h183;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h184;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h185;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h186;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h187;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h188;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h189;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h18f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h190;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h191;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h192;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h193;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h194;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h195;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h196;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h197;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h198;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h199;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h19f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h1ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h200;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h201;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h202;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h203;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h204;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h205;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h206;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h207;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h208;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h209;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h20f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h210;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h211;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h212;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h213;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h214;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h215;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h216;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h217;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h218;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h219;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h21f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h220;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h221;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h222;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h223;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h224;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h225;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h226;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h227;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h228;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h229;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h22f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h230;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h231;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h232;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h233;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h234;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h235;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h236;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h237;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h238;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h239;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h23f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h240;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h241;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h242;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h243;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h244;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h245;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h246;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h247;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h248;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h249;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h24f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h250;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h251;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h252;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h253;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h254;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h255;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h256;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h257;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h258;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h259;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h25f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h260;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h261;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h262;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h263;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h264;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h265;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h266;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h267;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h268;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h269;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h26f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h270;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h271;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h272;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h273;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h274;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h275;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h276;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h277;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h278;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h279;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h27f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h280;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h281;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h282;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h283;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h284;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h285;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h286;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h287;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h288;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h289;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h28f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h290;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h291;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h292;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h293;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h294;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h295;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h296;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h297;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h298;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h299;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h29f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h2ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h300;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h301;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h302;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h303;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h304;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h305;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h306;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h307;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h308;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h309;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h30f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h310;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h311;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h312;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h313;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h314;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h315;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h316;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h317;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h318;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h319;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h31f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h320;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h321;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h322;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h323;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h324;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h325;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h326;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h327;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h328;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h329;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h32f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h330;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h331;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h332;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h333;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h334;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h335;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h336;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h337;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h338;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h339;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h33f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h340;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h341;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h342;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h343;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h344;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h345;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h346;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h347;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h348;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h349;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h34f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h350;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h351;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h352;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h353;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h354;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h355;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h356;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h357;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h358;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h359;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h35f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h360;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h361;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h362;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h363;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h364;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h365;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h366;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h367;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h368;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h369;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h36f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h370;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h371;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h372;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h373;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h374;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h375;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h376;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h377;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h378;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h379;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h37f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h380;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h381;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h382;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h383;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h384;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h385;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h386;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h387;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h388;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h389;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h38f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h390;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h391;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h392;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h393;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h394;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h395;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h396;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h397;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h398;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h399;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h39f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h3ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h400;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h401;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h402;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h403;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h404;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h405;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h406;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h407;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h408;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h409;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h40f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h410;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h411;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h412;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h413;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h414;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h415;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h416;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h417;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h418;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h419;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h41f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h420;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h421;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h422;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h423;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h424;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h425;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h426;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h427;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h428;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h429;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h42f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h430;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h431;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h432;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h433;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h434;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h435;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h436;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h437;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h438;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h439;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h43f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h440;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h441;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h442;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h443;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h444;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h445;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h446;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h447;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h448;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h449;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h44f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h450;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h451;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h452;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h453;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h454;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h455;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h456;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h457;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h458;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h459;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h45f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h460;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h461;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h462;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h463;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h464;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h465;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h466;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h467;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h468;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h469;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h46f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h470;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h471;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h472;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h473;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h474;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h475;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h476;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h477;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h478;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h479;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h47f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h480;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h481;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h482;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h483;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h484;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h485;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h486;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h487;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h488;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h489;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h48f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h490;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h491;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h492;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h493;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h494;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h495;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h496;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h497;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h498;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h499;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h49f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h4ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h500;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h501;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h502;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h503;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h504;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h505;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h506;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h507;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h508;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h509;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h50f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h510;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h511;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h512;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h513;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h514;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h515;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h516;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h517;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h518;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h519;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h51f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h520;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h521;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h522;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h523;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h524;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h525;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h526;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h527;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h528;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h529;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h52f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h530;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h531;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h532;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h533;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h534;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h535;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h536;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h537;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h538;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h539;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h53f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h540;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h541;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h542;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h543;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h544;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h545;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h546;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h547;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h548;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h549;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h54f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h550;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h551;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h552;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h553;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h554;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h555;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h556;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h557;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h558;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h559;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h55f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h560;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h561;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h562;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h563;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h564;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h565;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h566;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h567;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h568;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h569;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h56f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h570;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h571;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h572;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h573;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h574;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h575;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h576;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h577;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h578;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h579;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h57f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h580;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h581;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h582;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h583;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h584;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h585;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h586;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h587;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h588;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h589;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h58f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h590;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h591;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h592;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h593;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h594;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h595;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h596;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h597;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h598;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h599;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h59f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h5ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h600;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h601;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h602;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h603;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h604;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h605;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h606;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h607;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h608;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h609;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h60f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h610;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h611;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h612;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h613;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h614;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h615;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h616;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h617;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h618;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h619;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h61f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h620;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h621;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h622;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h623;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h624;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h625;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h626;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h627;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h628;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h629;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h62f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h630;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h631;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h632;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h633;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h634;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h635;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h636;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h637;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h638;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h639;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h63f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h640;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h641;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h642;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h643;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h644;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h645;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h646;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h647;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h648;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h649;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h64f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h650;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h651;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h652;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h653;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h654;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h655;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h656;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h657;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h658;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h659;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h65f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h660;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h661;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h662;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h663;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h664;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h665;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h666;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h667;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h668;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h669;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h66f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h670;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h671;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h672;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h673;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h674;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h675;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h676;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h677;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h678;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h679;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h67f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h680;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h681;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h682;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h683;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h684;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h685;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h686;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h687;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h688;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h689;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h68f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h690;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h691;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h692;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h693;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h694;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h695;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h696;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h697;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h698;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h699;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h69f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h6ff;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h700;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h701;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h702;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h703;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h704;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h705;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h706;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h707;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h708;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h709;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h70f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h710;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h711;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h712;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h713;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h714;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h715;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h716;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h717;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h718;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h719;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h71f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h720;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h721;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h722;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h723;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h724;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h725;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h726;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h727;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h728;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h729;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h72f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h730;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h731;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h732;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h733;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h734;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h735;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h736;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h737;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h738;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h739;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h73f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h740;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h741;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h742;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h743;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h744;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h745;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h746;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h747;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h748;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h749;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h74f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h750;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h751;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h752;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h753;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h754;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h755;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h756;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h757;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h758;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h759;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h75f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h760;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h761;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h762;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h763;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h764;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h765;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h766;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h767;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h768;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h769;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h76f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h770;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h771;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h772;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h773;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h774;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h775;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h776;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h777;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h778;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h779;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h77f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h780;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h781;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h782;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h783;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h784;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h785;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h786;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h787;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h788;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h789;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h78f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h790;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h791;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h792;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h793;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h794;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h795;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h796;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h797;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h798;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h799;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79a;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79b;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79c;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79d;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79e;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h79f;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7a9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7aa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ab;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ac;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ad;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ae;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7af;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7b9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ba;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7bb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7bc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7bd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7be;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7bf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7c9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ca;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7cb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7cc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7cd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ce;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7cf;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7d9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7da;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7db;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7dc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7dd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7de;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7df;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7e9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ea;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7eb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ec;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ed;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ee;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ef;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f0;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f1;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f2;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f3;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f4;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f5;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f6;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f7;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f8;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7f9;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7fa;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7fb;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7fc;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7fd;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7fe;
        #1
        {src3[0], src2[3], src2[2], src2[1], src2[0], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 11'h7ff;
        #1
        $finish();
    end
endmodule
