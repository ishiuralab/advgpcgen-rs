module testbench();
    reg [4:0] src0;
    reg [2:0] src1;
    reg [0:0] src2;
    wire [3:0] dst;
    wire [3:0] exp;
    wire test;
    gpc135_4 gpc135_4(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .dst(dst)
    );
    assign exp = src0[0] * 1 + src0[1] * 1 + src0[2] * 1 + src0[3] * 1 + src0[4] * 1 + src1[0] * 2 + src1[1] * 2 + src1[2] * 2 + src2[0] * 4;
    assign test = dst == exp;
    initial begin
        $monitor("src0:0x%x, src1:0x%x, src2:0x%x, dst:0x%x, exp:0x%x, test:%x", src0, src1, src2, dst, exp, test);
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h20;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h21;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h22;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h23;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h24;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h25;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h26;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h27;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h28;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h29;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h2f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h30;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h31;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h32;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h33;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h34;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h35;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h36;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h37;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h38;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h39;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h3f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h40;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h41;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h42;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h43;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h44;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h45;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h46;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h47;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h48;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h49;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h4f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h50;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h51;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h52;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h53;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h54;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h55;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h56;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h57;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h58;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h59;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h5f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h60;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h61;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h62;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h63;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h64;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h65;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h66;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h67;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h68;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h69;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h6f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h70;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h71;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h72;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h73;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h74;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h75;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h76;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h77;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h78;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h79;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h7f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h80;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h81;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h82;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h83;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h84;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h85;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h86;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h87;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h88;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h89;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h8f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h90;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h91;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h92;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h93;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h94;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h95;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h96;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h97;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h98;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h99;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h9f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'ha9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'haa;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hab;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hac;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'had;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hae;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'haf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hb9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hba;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hbb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hbc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hbd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hbe;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hbf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hc9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hca;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hcb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hcc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hcd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hce;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hcf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hd9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hda;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hdb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hdc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hdd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hde;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hdf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'he9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hea;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'heb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hec;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hed;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hee;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hef;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hf9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hfa;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hfb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hfc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hfd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hfe;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'hff;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h100;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h101;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h102;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h103;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h104;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h105;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h106;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h107;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h108;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h109;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h10f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h110;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h111;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h112;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h113;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h114;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h115;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h116;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h117;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h118;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h119;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h11f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h120;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h121;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h122;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h123;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h124;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h125;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h126;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h127;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h128;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h129;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h12f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h130;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h131;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h132;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h133;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h134;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h135;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h136;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h137;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h138;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h139;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h13f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h140;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h141;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h142;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h143;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h144;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h145;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h146;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h147;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h148;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h149;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h14f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h150;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h151;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h152;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h153;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h154;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h155;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h156;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h157;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h158;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h159;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h15f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h160;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h161;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h162;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h163;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h164;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h165;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h166;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h167;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h168;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h169;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h16f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h170;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h171;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h172;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h173;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h174;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h175;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h176;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h177;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h178;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h179;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h17f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h180;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h181;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h182;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h183;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h184;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h185;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h186;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h187;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h188;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h189;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h18f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h190;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h191;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h192;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h193;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h194;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h195;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h196;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h197;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h198;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h199;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19a;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19b;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19c;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19d;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19e;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h19f;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1a9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1aa;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ab;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ac;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ad;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ae;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1af;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1b9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ba;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1bb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1bc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1bd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1be;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1bf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1c9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ca;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1cb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1cc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1cd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ce;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1cf;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1d9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1da;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1db;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1dc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1dd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1de;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1df;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1e9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ea;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1eb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ec;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ed;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ee;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ef;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f0;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f1;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f2;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f3;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f4;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f5;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f6;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f7;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f8;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1f9;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1fa;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1fb;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1fc;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1fd;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1fe;
        #1
        {src2[0], src1[2], src1[1], src1[0], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 9'h1ff;
        #1
        $finish();
    end
endmodule
