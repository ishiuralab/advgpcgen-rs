module testbench();
    reg [6:0] src0;
    reg [5:0] src2;
    wire [4:0] dst;
    wire [4:0] exp;
    wire test;
    gpc607_5 gpc607_5(
        .src0(src0),
        .src2(src2),
        .dst(dst)
    );
    assign exp = src0[0] * 1 + src0[1] * 1 + src0[2] * 1 + src0[3] * 1 + src0[4] * 1 + src0[5] * 1 + src0[6] * 1 + src2[0] * 4 + src2[1] * 4 + src2[2] * 4 + src2[3] * 4 + src2[4] * 4 + src2[5] * 4;
    assign test = dst == exp;
    initial begin
        $monitor("src0:0x%x, src2:0x%x, dst:0x%x, exp:0x%x, test:%x", src0, src2, dst, exp, test);
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h200;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h201;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h202;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h203;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h204;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h205;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h206;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h207;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h208;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h209;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h20f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h210;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h211;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h212;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h213;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h214;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h215;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h216;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h217;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h218;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h219;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h21f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h220;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h221;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h222;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h223;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h224;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h225;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h226;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h227;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h228;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h229;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h22f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h230;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h231;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h232;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h233;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h234;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h235;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h236;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h237;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h238;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h239;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h23f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h240;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h241;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h242;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h243;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h244;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h245;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h246;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h247;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h248;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h249;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h24f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h250;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h251;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h252;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h253;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h254;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h255;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h256;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h257;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h258;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h259;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h25f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h260;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h261;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h262;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h263;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h264;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h265;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h266;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h267;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h268;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h269;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h26f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h270;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h271;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h272;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h273;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h274;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h275;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h276;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h277;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h278;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h279;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h27f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h280;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h281;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h282;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h283;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h284;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h285;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h286;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h287;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h288;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h289;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h28f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h290;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h291;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h292;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h293;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h294;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h295;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h296;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h297;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h298;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h299;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h29f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h2ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h300;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h301;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h302;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h303;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h304;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h305;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h306;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h307;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h308;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h309;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h30f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h310;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h311;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h312;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h313;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h314;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h315;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h316;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h317;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h318;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h319;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h31f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h320;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h321;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h322;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h323;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h324;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h325;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h326;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h327;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h328;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h329;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h32f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h330;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h331;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h332;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h333;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h334;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h335;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h336;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h337;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h338;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h339;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h33f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h340;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h341;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h342;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h343;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h344;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h345;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h346;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h347;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h348;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h349;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h34f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h350;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h351;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h352;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h353;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h354;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h355;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h356;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h357;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h358;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h359;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h35f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h360;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h361;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h362;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h363;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h364;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h365;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h366;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h367;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h368;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h369;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h36f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h370;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h371;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h372;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h373;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h374;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h375;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h376;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h377;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h378;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h379;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h37f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h380;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h381;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h382;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h383;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h384;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h385;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h386;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h387;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h388;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h389;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h38f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h390;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h391;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h392;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h393;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h394;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h395;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h396;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h397;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h398;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h399;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h39f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h3ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h400;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h401;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h402;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h403;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h404;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h405;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h406;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h407;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h408;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h409;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h40f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h410;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h411;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h412;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h413;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h414;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h415;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h416;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h417;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h418;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h419;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h41f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h420;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h421;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h422;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h423;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h424;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h425;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h426;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h427;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h428;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h429;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h42f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h430;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h431;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h432;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h433;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h434;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h435;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h436;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h437;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h438;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h439;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h43f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h440;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h441;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h442;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h443;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h444;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h445;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h446;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h447;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h448;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h449;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h44f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h450;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h451;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h452;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h453;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h454;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h455;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h456;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h457;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h458;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h459;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h45f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h460;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h461;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h462;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h463;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h464;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h465;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h466;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h467;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h468;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h469;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h46f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h470;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h471;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h472;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h473;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h474;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h475;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h476;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h477;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h478;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h479;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h47f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h480;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h481;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h482;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h483;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h484;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h485;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h486;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h487;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h488;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h489;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h48f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h490;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h491;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h492;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h493;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h494;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h495;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h496;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h497;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h498;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h499;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h49f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h4ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h500;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h501;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h502;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h503;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h504;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h505;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h506;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h507;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h508;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h509;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h50f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h510;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h511;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h512;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h513;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h514;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h515;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h516;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h517;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h518;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h519;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h51f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h520;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h521;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h522;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h523;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h524;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h525;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h526;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h527;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h528;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h529;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h52f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h530;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h531;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h532;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h533;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h534;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h535;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h536;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h537;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h538;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h539;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h53f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h540;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h541;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h542;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h543;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h544;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h545;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h546;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h547;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h548;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h549;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h54f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h550;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h551;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h552;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h553;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h554;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h555;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h556;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h557;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h558;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h559;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h55f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h560;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h561;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h562;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h563;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h564;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h565;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h566;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h567;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h568;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h569;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h56f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h570;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h571;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h572;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h573;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h574;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h575;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h576;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h577;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h578;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h579;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h57f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h580;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h581;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h582;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h583;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h584;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h585;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h586;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h587;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h588;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h589;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h58f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h590;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h591;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h592;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h593;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h594;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h595;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h596;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h597;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h598;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h599;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h59f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h5ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h600;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h601;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h602;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h603;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h604;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h605;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h606;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h607;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h608;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h609;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h60f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h610;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h611;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h612;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h613;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h614;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h615;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h616;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h617;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h618;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h619;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h61f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h620;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h621;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h622;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h623;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h624;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h625;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h626;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h627;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h628;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h629;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h62f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h630;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h631;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h632;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h633;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h634;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h635;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h636;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h637;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h638;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h639;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h63f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h640;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h641;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h642;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h643;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h644;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h645;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h646;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h647;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h648;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h649;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h64f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h650;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h651;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h652;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h653;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h654;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h655;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h656;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h657;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h658;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h659;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h65f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h660;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h661;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h662;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h663;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h664;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h665;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h666;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h667;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h668;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h669;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h66f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h670;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h671;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h672;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h673;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h674;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h675;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h676;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h677;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h678;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h679;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h67f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h680;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h681;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h682;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h683;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h684;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h685;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h686;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h687;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h688;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h689;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h68f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h690;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h691;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h692;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h693;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h694;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h695;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h696;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h697;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h698;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h699;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h69f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h6ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h700;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h701;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h702;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h703;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h704;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h705;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h706;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h707;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h708;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h709;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h70f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h710;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h711;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h712;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h713;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h714;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h715;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h716;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h717;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h718;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h719;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h71f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h720;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h721;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h722;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h723;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h724;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h725;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h726;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h727;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h728;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h729;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h72f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h730;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h731;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h732;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h733;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h734;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h735;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h736;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h737;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h738;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h739;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h73f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h740;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h741;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h742;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h743;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h744;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h745;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h746;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h747;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h748;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h749;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h74f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h750;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h751;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h752;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h753;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h754;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h755;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h756;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h757;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h758;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h759;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h75f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h760;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h761;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h762;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h763;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h764;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h765;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h766;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h767;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h768;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h769;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h76f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h770;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h771;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h772;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h773;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h774;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h775;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h776;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h777;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h778;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h779;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h77f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h780;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h781;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h782;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h783;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h784;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h785;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h786;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h787;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h788;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h789;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h78f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h790;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h791;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h792;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h793;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h794;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h795;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h796;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h797;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h798;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h799;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h79f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h7ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h800;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h801;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h802;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h803;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h804;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h805;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h806;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h807;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h808;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h809;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h80f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h810;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h811;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h812;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h813;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h814;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h815;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h816;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h817;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h818;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h819;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h81f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h820;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h821;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h822;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h823;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h824;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h825;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h826;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h827;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h828;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h829;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h82f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h830;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h831;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h832;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h833;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h834;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h835;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h836;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h837;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h838;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h839;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h83f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h840;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h841;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h842;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h843;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h844;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h845;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h846;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h847;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h848;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h849;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h84f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h850;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h851;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h852;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h853;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h854;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h855;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h856;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h857;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h858;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h859;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h85f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h860;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h861;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h862;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h863;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h864;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h865;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h866;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h867;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h868;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h869;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h86f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h870;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h871;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h872;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h873;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h874;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h875;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h876;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h877;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h878;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h879;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h87f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h880;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h881;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h882;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h883;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h884;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h885;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h886;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h887;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h888;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h889;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h88f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h890;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h891;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h892;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h893;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h894;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h895;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h896;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h897;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h898;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h899;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h89f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h8ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h900;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h901;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h902;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h903;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h904;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h905;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h906;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h907;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h908;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h909;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h90f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h910;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h911;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h912;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h913;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h914;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h915;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h916;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h917;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h918;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h919;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h91f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h920;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h921;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h922;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h923;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h924;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h925;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h926;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h927;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h928;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h929;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h92f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h930;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h931;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h932;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h933;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h934;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h935;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h936;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h937;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h938;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h939;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h93f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h940;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h941;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h942;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h943;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h944;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h945;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h946;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h947;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h948;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h949;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h94f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h950;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h951;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h952;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h953;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h954;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h955;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h956;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h957;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h958;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h959;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h95f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h960;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h961;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h962;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h963;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h964;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h965;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h966;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h967;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h968;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h969;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h96f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h970;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h971;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h972;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h973;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h974;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h975;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h976;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h977;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h978;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h979;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h97f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h980;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h981;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h982;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h983;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h984;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h985;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h986;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h987;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h988;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h989;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h98f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h990;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h991;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h992;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h993;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h994;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h995;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h996;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h997;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h998;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h999;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h99f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h9ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'ha9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haa9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hab9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'habb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'habc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'habd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'habe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'habf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hac9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hacb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hacc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hacd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hace;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hacf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'had9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hada;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hadb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hadc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hadd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hade;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hadf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hae9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hafa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hafb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hafc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hafd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hafe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'haff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hb9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hba9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbe9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hbff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hc9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hca9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hccb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hccc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hccd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hccf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hce9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hceb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hced;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hcff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hd9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hda9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hddb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hddc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hddd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hddf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hde9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hded;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hdff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'he9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hea9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'head;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hebb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hebc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hebd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hebe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hebf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hec9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hecb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hecc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hecd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hece;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hecf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hed9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hedb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hedc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hedd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hede;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hedf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hee9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hef9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hefa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hefb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hefc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hefd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hefe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'heff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hf9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfa9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfe9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hff9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hffa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hffb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hffc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hffd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hffe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'hfff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1000;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1001;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1002;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1003;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1004;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1005;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1006;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1007;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1008;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1009;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h100f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1010;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1011;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1012;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1013;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1014;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1015;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1016;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1017;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1018;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1019;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h101f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1020;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1021;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1022;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1023;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1024;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1025;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1026;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1027;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1028;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1029;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h102f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1030;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1031;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1032;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1033;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1034;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1035;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1036;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1037;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1038;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1039;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h103f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1040;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1041;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1042;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1043;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1044;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1045;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1046;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1047;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1048;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1049;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h104f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1050;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1051;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1052;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1053;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1054;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1055;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1056;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1057;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1058;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1059;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h105f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1060;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1061;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1062;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1063;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1064;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1065;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1066;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1067;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1068;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1069;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h106f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1070;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1071;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1072;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1073;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1074;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1075;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1076;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1077;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1078;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1079;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h107f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1080;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1081;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1082;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1083;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1084;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1085;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1086;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1087;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1088;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1089;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h108f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1090;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1091;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1092;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1093;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1094;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1095;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1096;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1097;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1098;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1099;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h109f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h10ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1100;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1101;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1102;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1103;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1104;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1105;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1106;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1107;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1108;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1109;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h110f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1110;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1111;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1112;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1113;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1114;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1115;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1116;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1117;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1118;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1119;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h111f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1120;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1121;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1122;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1123;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1124;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1125;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1126;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1127;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1128;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1129;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h112f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1130;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1131;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1132;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1133;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1134;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1135;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1136;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1137;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1138;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1139;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h113f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1140;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1141;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1142;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1143;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1144;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1145;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1146;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1147;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1148;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1149;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h114f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1150;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1151;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1152;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1153;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1154;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1155;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1156;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1157;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1158;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1159;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h115f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1160;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1161;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1162;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1163;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1164;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1165;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1166;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1167;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1168;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1169;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h116f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1170;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1171;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1172;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1173;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1174;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1175;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1176;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1177;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1178;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1179;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h117f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1180;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1181;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1182;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1183;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1184;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1185;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1186;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1187;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1188;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1189;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h118f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1190;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1191;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1192;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1193;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1194;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1195;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1196;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1197;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1198;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1199;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h119f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h11ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1200;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1201;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1202;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1203;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1204;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1205;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1206;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1207;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1208;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1209;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h120f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1210;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1211;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1212;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1213;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1214;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1215;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1216;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1217;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1218;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1219;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h121f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1220;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1221;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1222;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1223;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1224;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1225;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1226;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1227;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1228;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1229;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h122f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1230;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1231;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1232;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1233;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1234;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1235;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1236;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1237;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1238;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1239;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h123f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1240;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1241;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1242;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1243;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1244;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1245;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1246;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1247;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1248;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1249;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h124f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1250;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1251;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1252;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1253;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1254;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1255;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1256;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1257;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1258;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1259;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h125f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1260;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1261;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1262;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1263;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1264;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1265;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1266;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1267;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1268;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1269;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h126f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1270;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1271;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1272;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1273;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1274;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1275;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1276;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1277;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1278;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1279;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h127f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1280;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1281;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1282;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1283;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1284;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1285;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1286;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1287;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1288;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1289;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h128f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1290;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1291;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1292;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1293;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1294;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1295;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1296;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1297;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1298;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1299;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h129f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h12ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1300;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1301;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1302;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1303;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1304;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1305;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1306;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1307;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1308;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1309;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h130f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1310;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1311;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1312;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1313;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1314;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1315;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1316;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1317;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1318;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1319;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h131f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1320;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1321;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1322;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1323;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1324;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1325;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1326;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1327;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1328;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1329;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h132f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1330;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1331;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1332;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1333;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1334;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1335;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1336;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1337;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1338;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1339;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h133f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1340;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1341;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1342;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1343;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1344;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1345;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1346;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1347;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1348;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1349;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h134f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1350;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1351;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1352;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1353;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1354;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1355;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1356;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1357;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1358;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1359;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h135f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1360;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1361;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1362;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1363;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1364;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1365;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1366;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1367;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1368;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1369;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h136f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1370;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1371;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1372;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1373;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1374;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1375;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1376;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1377;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1378;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1379;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h137f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1380;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1381;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1382;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1383;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1384;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1385;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1386;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1387;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1388;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1389;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h138f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1390;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1391;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1392;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1393;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1394;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1395;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1396;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1397;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1398;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1399;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h139f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h13ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1400;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1401;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1402;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1403;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1404;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1405;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1406;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1407;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1408;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1409;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h140f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1410;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1411;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1412;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1413;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1414;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1415;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1416;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1417;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1418;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1419;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h141f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1420;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1421;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1422;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1423;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1424;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1425;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1426;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1427;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1428;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1429;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h142f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1430;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1431;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1432;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1433;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1434;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1435;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1436;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1437;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1438;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1439;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h143f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1440;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1441;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1442;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1443;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1444;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1445;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1446;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1447;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1448;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1449;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h144f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1450;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1451;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1452;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1453;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1454;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1455;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1456;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1457;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1458;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1459;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h145f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1460;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1461;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1462;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1463;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1464;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1465;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1466;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1467;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1468;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1469;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h146f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1470;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1471;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1472;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1473;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1474;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1475;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1476;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1477;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1478;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1479;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h147f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1480;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1481;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1482;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1483;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1484;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1485;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1486;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1487;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1488;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1489;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h148f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1490;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1491;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1492;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1493;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1494;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1495;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1496;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1497;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1498;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1499;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h149f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h14ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1500;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1501;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1502;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1503;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1504;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1505;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1506;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1507;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1508;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1509;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h150f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1510;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1511;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1512;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1513;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1514;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1515;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1516;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1517;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1518;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1519;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h151f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1520;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1521;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1522;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1523;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1524;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1525;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1526;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1527;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1528;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1529;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h152f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1530;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1531;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1532;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1533;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1534;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1535;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1536;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1537;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1538;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1539;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h153f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1540;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1541;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1542;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1543;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1544;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1545;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1546;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1547;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1548;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1549;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h154f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1550;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1551;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1552;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1553;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1554;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1555;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1556;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1557;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1558;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1559;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h155f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1560;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1561;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1562;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1563;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1564;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1565;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1566;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1567;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1568;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1569;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h156f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1570;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1571;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1572;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1573;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1574;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1575;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1576;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1577;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1578;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1579;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h157f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1580;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1581;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1582;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1583;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1584;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1585;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1586;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1587;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1588;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1589;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h158f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1590;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1591;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1592;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1593;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1594;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1595;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1596;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1597;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1598;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1599;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h159f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h15ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1600;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1601;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1602;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1603;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1604;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1605;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1606;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1607;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1608;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1609;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h160f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1610;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1611;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1612;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1613;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1614;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1615;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1616;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1617;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1618;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1619;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h161f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1620;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1621;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1622;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1623;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1624;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1625;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1626;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1627;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1628;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1629;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h162f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1630;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1631;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1632;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1633;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1634;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1635;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1636;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1637;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1638;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1639;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h163f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1640;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1641;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1642;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1643;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1644;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1645;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1646;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1647;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1648;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1649;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h164f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1650;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1651;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1652;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1653;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1654;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1655;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1656;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1657;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1658;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1659;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h165f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1660;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1661;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1662;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1663;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1664;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1665;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1666;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1667;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1668;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1669;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h166f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1670;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1671;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1672;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1673;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1674;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1675;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1676;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1677;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1678;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1679;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h167f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1680;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1681;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1682;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1683;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1684;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1685;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1686;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1687;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1688;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1689;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h168f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1690;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1691;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1692;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1693;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1694;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1695;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1696;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1697;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1698;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1699;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h169f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h16ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1700;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1701;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1702;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1703;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1704;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1705;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1706;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1707;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1708;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1709;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h170f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1710;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1711;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1712;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1713;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1714;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1715;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1716;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1717;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1718;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1719;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h171f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1720;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1721;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1722;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1723;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1724;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1725;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1726;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1727;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1728;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1729;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h172f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1730;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1731;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1732;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1733;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1734;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1735;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1736;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1737;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1738;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1739;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h173f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1740;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1741;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1742;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1743;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1744;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1745;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1746;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1747;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1748;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1749;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h174f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1750;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1751;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1752;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1753;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1754;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1755;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1756;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1757;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1758;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1759;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h175f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1760;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1761;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1762;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1763;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1764;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1765;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1766;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1767;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1768;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1769;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h176f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1770;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1771;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1772;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1773;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1774;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1775;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1776;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1777;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1778;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1779;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h177f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1780;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1781;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1782;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1783;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1784;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1785;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1786;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1787;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1788;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1789;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h178f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1790;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1791;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1792;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1793;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1794;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1795;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1796;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1797;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1798;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1799;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h179f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h17ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1800;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1801;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1802;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1803;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1804;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1805;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1806;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1807;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1808;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1809;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h180f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1810;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1811;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1812;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1813;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1814;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1815;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1816;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1817;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1818;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1819;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h181f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1820;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1821;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1822;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1823;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1824;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1825;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1826;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1827;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1828;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1829;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h182f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1830;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1831;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1832;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1833;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1834;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1835;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1836;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1837;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1838;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1839;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h183f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1840;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1841;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1842;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1843;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1844;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1845;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1846;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1847;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1848;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1849;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h184f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1850;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1851;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1852;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1853;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1854;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1855;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1856;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1857;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1858;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1859;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h185f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1860;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1861;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1862;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1863;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1864;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1865;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1866;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1867;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1868;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1869;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h186f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1870;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1871;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1872;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1873;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1874;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1875;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1876;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1877;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1878;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1879;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h187f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1880;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1881;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1882;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1883;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1884;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1885;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1886;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1887;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1888;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1889;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h188f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1890;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1891;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1892;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1893;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1894;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1895;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1896;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1897;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1898;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1899;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h189f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h18ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1900;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1901;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1902;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1903;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1904;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1905;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1906;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1907;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1908;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1909;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h190f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1910;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1911;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1912;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1913;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1914;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1915;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1916;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1917;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1918;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1919;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h191f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1920;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1921;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1922;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1923;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1924;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1925;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1926;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1927;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1928;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1929;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h192f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1930;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1931;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1932;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1933;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1934;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1935;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1936;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1937;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1938;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1939;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h193f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1940;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1941;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1942;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1943;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1944;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1945;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1946;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1947;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1948;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1949;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h194f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1950;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1951;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1952;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1953;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1954;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1955;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1956;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1957;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1958;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1959;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h195f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1960;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1961;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1962;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1963;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1964;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1965;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1966;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1967;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1968;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1969;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h196f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1970;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1971;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1972;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1973;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1974;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1975;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1976;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1977;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1978;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1979;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h197f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1980;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1981;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1982;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1983;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1984;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1985;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1986;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1987;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1988;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1989;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h198f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1990;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1991;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1992;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1993;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1994;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1995;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1996;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1997;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1998;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1999;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h199f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19a9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19aa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19af;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19b9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19bb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19bc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19bd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19be;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19bf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19c9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19cb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19cc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19cd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19cf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19d9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19da;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19db;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19dc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19dd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19de;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19df;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19e9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19eb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19f9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19fa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19fb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19fc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19fd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19fe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h19ff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1a9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aa9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ab9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1abb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1abc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1abd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1abe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1abf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ac9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1acb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1acc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1acd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ace;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1acf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ad9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ada;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1adb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1adc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1add;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ade;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1adf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ae9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1af9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1afa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1afb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1afc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1afd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1afe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1aff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1b9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ba9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1baa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1baf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1be9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1beb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1bff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1c9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ca9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1caa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1caf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ccb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ccc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ccd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ccf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ce9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ceb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ced;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cf9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1cff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1d9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1da9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1daa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1daf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1db9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ddb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ddc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ddd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ddf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1de9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1deb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ded;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1def;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1df9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dfa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dfb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dfc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dfd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dfe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1dff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1e9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ea9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eaa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ead;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eaf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ebb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ebc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ebd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ebe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ebf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ec9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ecb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ecc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ecd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ece;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ecf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ed9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1edb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1edc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1edd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ede;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1edf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ee9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eeb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ef9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1efa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1efb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1efc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1efd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1efe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1eff;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f00;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f01;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f02;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f03;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f04;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f05;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f06;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f07;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f08;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f09;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f0f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f10;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f11;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f12;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f13;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f14;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f15;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f16;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f17;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f18;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f19;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f1f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f20;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f21;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f22;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f23;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f24;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f25;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f26;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f27;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f28;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f29;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f2f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f30;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f31;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f32;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f33;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f34;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f35;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f36;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f37;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f38;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f39;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f3f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f40;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f41;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f42;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f43;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f44;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f45;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f46;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f47;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f48;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f49;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f4f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f50;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f51;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f52;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f53;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f54;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f55;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f56;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f57;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f58;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f59;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f5f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f60;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f61;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f62;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f63;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f64;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f65;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f66;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f67;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f68;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f69;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f6f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f70;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f71;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f72;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f73;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f74;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f75;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f76;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f77;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f78;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f79;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f7f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f80;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f81;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f82;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f83;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f84;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f85;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f86;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f87;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f88;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f89;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f8f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f90;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f91;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f92;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f93;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f94;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f95;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f96;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f97;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f98;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f99;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9a;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9b;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9c;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9d;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9e;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1f9f;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fa9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1faa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fab;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fac;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fad;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fae;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1faf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fb9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fba;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fbb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fbc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fbd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fbe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fbf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fc9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fca;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fcb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fcc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fcd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fce;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fcf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fd9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fda;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fdb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fdc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fdd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fde;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fdf;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fe9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fea;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1feb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fec;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fed;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fee;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fef;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff0;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff1;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff2;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff3;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff4;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff5;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff6;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff7;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff8;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ff9;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ffa;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ffb;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ffc;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ffd;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1ffe;
        #1
        {src2[5], src2[4], src2[3], src2[2], src2[1], src2[0], src0[6], src0[5], src0[4], src0[3], src0[2], src0[1], src0[0]} <= 13'h1fff;
        #1
        $finish();
    end
endmodule
